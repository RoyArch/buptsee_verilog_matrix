module matrix(input wire clk,
		    		  input wire rst,
              output wire [7:0]col_r,
              output wire [7:0]col_g,
              output wire [7:0]row);
reg [63:0] temp;
reg[9:0]cnt;
reg[2:0]state;

matOut processer(
.char(temp),
.color(1'b0),
.clk(clk),
.rst(rst),
.row(row),
.col_r(col_r),
.col_g(col_g)
);

always@(posedge clk or posedge rst)
begin
  if(rst) begin
    cnt<=0;
    state<=0;
  end
  else begin
    if(cnt==10'd999)
    begin
      if(state>=3'd5) state<=3'd0;
      else state<=state+3'd1;
      cnt<=10'b0;
    end
	 else cnt<=cnt+10'b1;
  end
end

always@(*)
begin
  case(state)
  3'd0:temp=char_B;
  3'd1:temp=char_U;
  3'd2:temp=char_P;
  3'd3:temp=char_T;
  3'd4:temp=char_D;
  3'd5:temp=char_Y;
  endcase
end

parameter RED=0;
parameter GREEN=1;

parameter char_0 =64'h003C4242C2423C00;//0

parameter char_1 =64'h0018381818181800;//1

parameter char_2 =64'h003C460418207E00;//2

parameter char_3 =64'h003C460C16423C00;//3

parameter char_4 =64'h000C1C2C4CFE0C00;//4

parameter char_5 =64'h007E60FC02463C00;//5

parameter char_6 =64'h003E605C62623C00;//6

parameter char_7 =64'h007E040408081000;//7

parameter char_8 =64'h003C46245E423C00;//8

parameter char_9 =64'h003C46463A067800;//9

parameter char_A =64'h00181824247EC300;//A0

parameter char_B =64'h00FEC2FCC2C2FC00;//B1

parameter char_C =64'h003E424040433C00;//C2

parameter char_D =64'h00FCC2C2C2C6FC00;//D3

parameter char_E =64'h00FEC0FEC0C0FE00;//E4

parameter char_F =64'h00FEC0FCC0C0C000;//F5

parameter char_G =64'h003E42404E463E00;//G6

parameter char_H =64'h00C6C6FEC6C6C600;//H7

parameter char_I =64'h0018181818181800;//I8

parameter char_J =64'h00060606C6C63C00;//J9

parameter char_K =64'h00C6D8F0C8C4C700;//K10

parameter char_L =64'h00C0C0C0C0C0FE00;//L11

parameter char_M =64'h00C366665A52D700;//M12

parameter char_N =64'h00E6F6D6CECEC600;//N13

parameter char_O =64'h007C4242C2423C00;//O14

parameter char_P =64'h00FEC2C6FCC0C000;//P15

parameter char_Q =64'h007C4242C24E3E00;//Q16

parameter char_R =64'h00FEC2CEFCC4C700;//R17

parameter char_S =64'h003E42300E423C00;//S18

parameter char_T =64'h007E181818181800;//T19

parameter char_U =64'h00C6C6C6C6C67C00;//U20

parameter char_V =64'h00C366242C381800;//V21

parameter char_W =64'h00DBDA5A6E666600;//W22

parameter char_X =64'h00662C181824C700;//X23

parameter char_Y =64'h00C3243818181800;//Y24

parameter char_Z =64'h007E040810207E00;//Z25
endmodule